//: version "1.8.7"

module ALU_PLUS_MINUS(i22, i21, i12, o6, s, o12, i11, co);
//: interface  /sz:(40, 40) /bd:[ ]
input i11;    //: /sn:0 /dp:1 {0}(322,143)(42,143)(42,248)(-29,248){1}
input i21;    //: /sn:0 /dp:1 {0}(324,317)(68,317)(68,301)(-30,301){1}
output o12;    //: /sn:0 {0}(1715,308)(1572,308)(1572,320)(1556,320){1}
input i12;    //: /sn:0 /dp:1 {0}(318,233)(81,233)(81,273)(-31,273){1}
output co;    //: /sn:0 {0}(1715,327)(1619,327)(1619,495)(1381,495){1}
input i22;    //: /sn:0 /dp:1 {0}(331,428)(39,428)(39,334)(-33,334){1}
input s;    //: /sn:0 /dp:13 {0}(1513,385)(1513,616)(1411,616){1}
//: {2}(1409,614)(1409,607)(1418,607)(1418,182){3}
//: {4}(1407,616)(1295,616){5}
//: {6}(1293,614)(1293,588)(1335,588)(1335,560){7}
//: {8}(1291,616)(382,616)(382,573)(226,573){9}
//: {10}(224,571)(224,423){11}
//: {12}(226,421)(248,421)(248,450)(331,450){13}
//: {14}(224,419)(224,349)(232,349){15}
//: {16}(236,349)(276,349){17}
//: {18}(280,349)(295,349)(295,339)(324,339){19}
//: {20}(278,347)(278,165)(322,165){21}
//: {22}(234,347)(234,255)(318,255){23}
//: {24}(222,573)(-6,573)(-6,353)(-33,353){25}
output o6;    //: /sn:0 {0}(1713,287)(1579,287)(1579,117)(1464,117){1}
wire w6;    //: /sn:0 {0}(429,317)(549,317)(549,276)(712,276){1}
wire o8;    //: /sn:0 {0}(423,261)(599,261)(599,490)(692,490){1}
wire o11;    //: /sn:0 {0}(436,456)(573,456)(573,554)(692,554){1}
wire co0;    //: /sn:0 {0}(1300,476)(1206,476)(1206,274)(901,274){1}
wire w3;    //: /sn:0 {0}(423,233)(653,233)(653,195)(712,195){1}
wire o1;    //: /sn:0 {0}(884,471)(1001,471)(1001,146)(1383,146){1}
wire o9;    //: /sn:0 {0}(884,492)(1149,492)(1149,349)(1475,349){1}
wire o7;    //: /sn:0 {0}(427,171)(633,171)(633,469)(692,469){1}
wire o3;    //: /sn:0 {0}(901,234)(1447,234)(1447,301)(1475,301){1}
wire w2;    //: /sn:0 {0}(427,143)(656,143)(656,180)(712,180){1}
wire o10;    //: /sn:0 {0}(429,345)(584,345)(584,536)(692,536){1}
wire i4;    //: /sn:0 {0}(1300,524)(973,524)(973,545)(884,545){1}
wire o2;    //: /sn:0 {0}(901,210)(1239,210)(1239,98)(1383,98){1}
wire w9;    //: /sn:0 {0}(436,428)(673,428)(673,294)(712,294){1}
//: enddecls

  //: input g4 (i22) @(-35,334) /sn:0 /w:[ 1 ]
  DEMUX g8 (.s(s), .i1(i12), .o2(o8), .o1(w3));   //: @(319, 210) /sz:(103, 75) /sn:0 /p:[ Li0>23 Li1>0 Ro0<0 Ro1<0 ]
  two_bit_FA g3 (.i22(w9), .i21(w6), .i12(w3), .i11(w2), .co(co0), .o2(o3), .o1(o2));   //: @(713, 147) /sz:(187, 190) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Ro0<1 Ro1<0 Ro2<0 ]
  DEMUX g13 (.s(s), .i1(i22), .o2(o11), .o1(w9));   //: @(332, 405) /sz:(103, 75) /sn:0 /p:[ Li0>13 Li1>0 Ro0<0 Ro1<0 ]
  //: input g2 (i21) @(-32,301) /sn:0 /w:[ 1 ]
  //: input g1 (i12) @(-33,273) /sn:0 /w:[ 1 ]
  //: joint g11 (s) @(224, 421) /w:[ 12 14 -1 11 ]
  //: joint g16 (s) @(1293, 616) /w:[ 5 6 8 -1 ]
  //: joint g10 (s) @(224, 573) /w:[ 9 10 24 -1 ]
  MUX g19 (.i2(co0), .i1(i4), .s(s), .o(co));   //: @(1301, 439) /sz:(79, 121) /sn:0 /p:[ Li0>0 Li1>0 Bi0>7 Ro0<1 ]
  DEMUX g6 (.s(s), .i1(i11), .o2(o7), .o1(w2));   //: @(323, 120) /sz:(103, 75) /sn:0 /p:[ Li0>21 Li1>0 Ro0<0 Ro1<0 ]
  //: joint g7 (s) @(234, 349) /w:[ 16 22 15 -1 ]
  //: joint g9 (s) @(278, 349) /w:[ 18 20 17 -1 ]
  MUX g15 (.i2(o2), .i1(o1), .s(s), .o(o6));   //: @(1384, 61) /sz:(79, 121) /sn:0 /p:[ Li0>1 Li1>1 Bi0>3 Ro0<1 ]
  //: output g20 (o6) @(1710,287) /sn:0 /w:[ 0 ]
  MUX g17 (.i2(o3), .i1(o9), .s(s), .o(o12));   //: @(1476, 264) /sz:(79, 121) /sn:0 /p:[ Li0>1 Li1>1 Bi0>0 Ro0<1 ]
  //: input g5 (s) @(-35,353) /sn:0 /w:[ 25 ]
  two_bit_sustractor g14 (.i22(o11), .i21(o10), .i12(o8), .i11(o7), .co(i4), .o2(o9), .o1(o1));   //: @(693, 422) /sz:(190, 162) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Ro0<1 Ro1<0 Ro2<0 ]
  //: output g21 (o12) @(1712,308) /sn:0 /w:[ 0 ]
  //: input g0 (i11) @(-31,248) /sn:0 /w:[ 1 ]
  //: output g22 (co) @(1712,327) /sn:0 /w:[ 0 ]
  DEMUX g12 (.s(s), .i1(i21), .o2(o10), .o1(w6));   //: @(325, 294) /sz:(103, 75) /sn:0 /p:[ Li0>19 Li1>0 Ro0<0 Ro1<0 ]
  //: joint g18 (s) @(1409, 616) /w:[ 1 2 4 -1 ]

endmodule

module MUX(i2, i1, o, s);
//: interface  /sz:(40, 40) /bd:[ ]
input i2;    //: /sn:0 /dp:1 {0}(365,309)(355,309)(355,294)(417,294)(417,203){1}
input i1;    //: /sn:0 {0}(332,207)(332,363)(365,363){1}
output o;    //: /sn:0 /dp:1 {0}(469,319)(552,319){1}
input s;    //: /sn:0 /dp:1 {0}(365,314)(177,314)(177,259){1}
//: {2}(179,257)(224,257)(224,334)(245,334){3}
//: {4}(175,257)(163,257){5}
wire w3;    //: /sn:0 /dp:1 {0}(448,321)(396,321)(396,366)(386,366){1}
wire w0;    //: /sn:0 /dp:1 {0}(448,316)(396,316)(396,312)(386,312){1}
wire w1;    //: /sn:0 /dp:1 {0}(365,368)(288,368)(288,334)(261,334){1}
//: enddecls

  or g8 (.I0(w0), .I1(w3), .Z(o));   //: @(459,319) /sn:0 /w:[ 0 0 0 ]
  not g4 (.I(s), .Z(w1));   //: @(251,334) /sn:0 /w:[ 3 1 ]
  and g3 (.I0(i2), .I1(s), .Z(w0));   //: @(376,312) /sn:0 /w:[ 0 0 1 ]
  //: input g2 (i2) @(417,201) /sn:0 /R:3 /w:[ 1 ]
  //: input g1 (i1) @(332,205) /sn:0 /R:3 /w:[ 0 ]
  and g6 (.I0(i1), .I1(w1), .Z(w3));   //: @(376,366) /sn:0 /w:[ 1 0 1 ]
  //: output g9 (o) @(549,319) /sn:0 /w:[ 1 ]
  //: joint g5 (s) @(177, 257) /w:[ 2 -1 4 1 ]
  //: input g0 (s) @(161,257) /sn:0 /w:[ 5 ]

endmodule

module HA(b, a, o, co);
//: interface  /sz:(40, 40) /bd:[ ]
input b;    //: /sn:0 {0}(433,306)(446,306){1}
//: {2}(450,306)(482,306)(482,284)(490,284){3}
//: {4}(448,308)(448,331)(503,331){5}
output co;    //: /sn:0 /dp:1 {0}(511,282)(596,282)(596,306)(606,306){1}
output o;    //: /sn:0 {0}(607,319)(579,319)(579,329)(524,329){1}
input a;    //: /sn:0 {0}(430,265)(466,265){1}
//: {2}(470,265)(482,265)(482,279)(490,279){3}
//: {4}(468,267)(468,326)(503,326){5}
//: enddecls

  //: joint g4 (a) @(468, 265) /w:[ 2 -1 1 4 ]
  //: input g3 (b) @(431,306) /sn:0 /w:[ 0 ]
  //: input g2 (a) @(428,265) /sn:0 /w:[ 0 ]
  xor g1 (.I0(a), .I1(b), .Z(o));   //: @(514,329) /sn:0 /w:[ 5 5 1 ]
  //: output g6 (o) @(604,319) /sn:0 /w:[ 0 ]
  //: output g7 (co) @(603,306) /sn:0 /w:[ 1 ]
  //: joint g5 (b) @(448, 306) /w:[ 2 -1 1 4 ]
  and g0 (.I0(a), .I1(b), .Z(co));   //: @(501,282) /sn:0 /w:[ 3 3 0 ]

endmodule

module two_bit_sustractor(i21, o1, i12, co, o2, i22, i11);
//: interface  /sz:(40, 40) /bd:[ ]
input i11;    //: /sn:0 {0}(76,195)(476,195)(476,202)(603,202){1}
input i21;    //: /sn:0 /dp:1 {0}(371,294)(260,294)(260,295)(78,295){1}
output o1;    //: /sn:0 {0}(982,232)(792,232){1}
input i12;    //: /sn:0 {0}(79,255)(80,255)(80,256)(127,256){1}
//: {2}(129,254)(129,217)(603,217){3}
//: {4}(129,258)(129,261){5}
output co;    //: /sn:0 {0}(986,274)(976,274)(976,314)(792,314){1}
input i22;    //: /sn:0 {0}(78,334)(261,334){1}
//: {2}(265,334)(595,334)(595,316)(603,316){3}
//: {4}(263,332)(263,299)(371,299){5}
output o2;    //: /sn:0 {0}(792,256)(974,256)(974,251)(984,251){1}
wire w3;    //: /sn:0 {0}(392,297)(533,297)(533,298)(603,298){1}
//: enddecls

  //: input g4 (i21) @(76,295) /sn:0 /w:[ 1 ]
  //: output g8 (o1) @(979,232) /sn:0 /w:[ 0 ]
  two_bit_FA g3 (.i22(i22), .i21(w3), .i12(i12), .i11(i11), .co(co), .o2(o2), .o1(o1));   //: @(604, 169) /sz:(187, 190) /sn:0 /p:[ Li0>3 Li1>1 Li2>3 Li3>1 Ro0<1 Ro1<0 Ro2<1 ]
  //: joint g2 (i12) @(129, 256) /w:[ -1 2 1 4 ]
  //: input g1 (i12) @(77,255) /sn:0 /w:[ 0 ]
  //: output g10 (co) @(983,274) /sn:0 /w:[ 0 ]
  xor g6 (.I0(i21), .I1(i22), .Z(w3));   //: @(382,297) /sn:0 /w:[ 0 5 0 ]
  //: joint g7 (i22) @(263, 334) /w:[ 2 4 1 -1 ]
  //: output g9 (o2) @(981,251) /sn:0 /w:[ 1 ]
  //: input g5 (i22) @(76,334) /sn:0 /w:[ 0 ]
  //: input g0 (i11) @(74,195) /sn:0 /w:[ 0 ]

endmodule

module DEMUX(o2, o1, s, i1);
//: interface  /sz:(40, 40) /bd:[ ]
output o1;    //: /sn:0 {0}(699,286)(688,286)(688,252)(530,252){1}
input i1;    //: /sn:0 {0}(168,284)(285,284){1}
//: {2}(289,284)(299,284)(299,298)(307,298){3}
//: {4}(287,282)(287,249)(509,249){5}
input s;    //: /sn:0 {0}(164,336)(286,336){1}
//: {2}(290,336)(299,336)(299,303)(307,303){3}
//: {4}(288,338)(288,363)(343,363){5}
output o2;    //: /sn:0 /dp:1 {0}(328,301)(555,301)(555,309)(700,309){1}
wire w1;    //: /sn:0 {0}(359,363)(433,363)(433,254)(509,254){1}
//: enddecls

  and g4 (.I0(i1), .I1(s), .Z(o2));   //: @(318,301) /sn:0 /w:[ 3 3 0 ]
  and g8 (.I0(i1), .I1(w1), .Z(o1));   //: @(520,252) /sn:0 /w:[ 5 1 1 ]
  //: output g3 (o2) @(697,309) /sn:0 /w:[ 1 ]
  //: output g2 (o1) @(696,286) /sn:0 /w:[ 0 ]
  //: input g1 (s) @(162,336) /sn:0 /w:[ 0 ]
  not g6 (.I(s), .Z(w1));   //: @(349,363) /sn:0 /w:[ 5 0 ]
  //: joint g7 (s) @(288, 336) /w:[ 2 -1 1 4 ]
  //: joint g9 (i1) @(287, 284) /w:[ 2 4 1 -1 ]
  //: input g0 (i1) @(166,284) /sn:0 /w:[ 0 ]

endmodule

module D2_bit_FA(i22, co, i21, i12, i11, o1, o2);
//: interface  /sz:(40, 40) /bd:[ ]
input i11;    //: /sn:0 {0}(635,152)(73,152)(73,221)(61,221){1}
input i21;    //: /sn:0 /dp:1 {0}(635,170)(358,170)(358,197)(108,197)(108,304)(67,304){1}
output o1;    //: /sn:0 {0}(922,340)(905,340)(905,385)(528,385){1}
input i12;    //: /sn:0 {0}(65,245)(325,245)(325,394)(386,394){1}
output co;    //: /sn:0 {0}(707,177)(912,177)(912,305)(922,305){1}
input i22;    //: /sn:0 {0}(67,335)(296,335)(296,442)(386,442){1}
output o2;    //: /sn:0 {0}(707,153)(851,153)(851,322)(922,322){1}
wire co0;    //: /sn:0 {0}(528,446)(625,446)(625,197)(635,197){1}
//: enddecls

  //: input g4 (i22) @(65,335) /sn:0 /w:[ 0 ]
  //: output g8 (co) @(919,305) /sn:0 /w:[ 1 ]
  //: input g3 (i21) @(65,304) /sn:0 /w:[ 1 ]
  //: input g2 (i12) @(63,245) /sn:0 /w:[ 0 ]
  //: input g1 (i11) @(59,221) /sn:0 /w:[ 1 ]
  HA g6 (.b(i22), .a(i12), .co(co0), .o(o1));   //: @(387, 346) /sz:(140, 123) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  //: output g7 (o1) @(919,340) /sn:0 /w:[ 0 ]
  FA g5 (.ci(co0), .b(i21), .a(i11), .co(co), .o(o2));   //: @(636, 131) /sz:(70, 92) /sn:0 /p:[ Li0>1 Li1>0 Li2>0 Ro0<0 Ro1<0 ]
  //: output g0 (o2) @(919,322) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(314,308)(446,308)(446,297)(456,297){1}
wire w7;    //: /sn:0 {0}(318,344)(446,344)(446,319)(456,319){1}
wire w4;    //: /sn:0 {0}(318,234)(437,234)(437,225)(456,225){1}
wire w3;    //: /sn:0 {0}(319,197)(408,197)(408,199)(456,199){1}
wire o12;    //: /sn:0 {0}(636,249)(626,249){1}
wire co2;    //: /sn:0 {0}(636,276)(626,276){1}
wire w5;    //: /sn:0 {0}(318,269)(446,269)(446,261)(456,261){1}
wire o6;    //: /sn:0 {0}(636,207)(626,207){1}
//: enddecls

  ALU_PLUS_MINUS g4 (.s(w7), .i22(w6), .i21(w5), .i12(w4), .i11(w3), .co(co2), .o12(o12), .o6(o6));   //: @(457, 151) /sz:(168, 192) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Ro0<1 Ro1<1 Ro2<1 ]
  //: switch g8 (w4) @(301,234) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w3) @(302,197) /sn:0 /w:[ 0 ] /st:1
  //: switch g11 (w7) @(301,344) /sn:0 /w:[ 0 ] /st:1
  //: switch g10 (w6) @(297,308) /sn:0 /w:[ 0 ] /st:1
  //: switch g9 (w5) @(301,269) /sn:0 /w:[ 0 ] /st:0

endmodule

module FA(ci, b, a, co, o);
//: interface  /sz:(40, 40) /bd:[ ]
input b;    //: /sn:0 {0}(-183,214)(95,214)(95,240)(103,240){1}
output co;    //: /sn:0 /dp:1 {0}(493,256)(756,256)(756,210)(766,210){1}
output o;    //: /sn:0 /dp:1 {0}(647,124)(755,124)(755,196)(765,196){1}
input ci;    //: /sn:0 {0}(-181,270)(341,270)(341,251)(351,251){1}
input a;    //: /sn:0 {0}(-178,133)(93,133)(93,192)(103,192){1}
wire co0;    //: /sn:0 {0}(245,244)(341,244)(341,195)(351,195){1}
wire w0;    //: /sn:0 {0}(493,184)(589,184)(589,126)(626,126){1}
wire o0;    //: /sn:0 {0}(245,183)(333,183)(333,121)(626,121){1}
//: enddecls

  //: input g4 (ci) @(-183,270) /sn:0 /w:[ 0 ]
  HA g3 (.b(ci), .a(co0), .co(co), .o(w0));   //: @(352, 139) /sz:(140, 144) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: input g2 (b) @(-185,214) /sn:0 /w:[ 0 ]
  //: input g1 (a) @(-180,133) /sn:0 /w:[ 0 ]
  //: output g6 (co) @(763,210) /sn:0 /w:[ 1 ]
  //: output g7 (o) @(762,196) /sn:0 /w:[ 1 ]
  or g5 (.I0(o0), .I1(w0), .Z(o));   //: @(637,124) /sn:0 /w:[ 1 1 0 ]
  HA g0 (.b(b), .a(a), .co(co0), .o(o0));   //: @(104, 144) /sz:(140, 123) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]

endmodule

module two_bit_FA(co, i22, i21, i12, o1, o2, i11);
//: interface  /sz:(40, 40) /bd:[ ]
input i11;    //: /sn:0 {0}(165,159)(550,159)(550,198)(560,198){1}
output o1;    //: /sn:0 {0}(856,214)(722,214)(722,200)(692,200){1}
input i21;    //: /sn:0 {0}(165,264)(460,264)(460,225)(560,225){1}
input i12;    //: /sn:0 {0}(165,184)(290,184)(290,328)(300,328){1}
output co;    //: /sn:0 {0}(858,237)(703,237)(703,235)(692,235){1}
input i22;    //: /sn:0 /dp:1 {0}(300,353)(174,353)(174,296)(166,296){1}
output o2;    //: /sn:0 {0}(405,327)(848,327)(848,259)(858,259){1}
wire co0;    //: /sn:0 {0}(405,349)(506,349)(506,246)(560,246){1}
//: enddecls

  //: output g8 (co) @(855,237) /sn:0 /w:[ 0 ]
  FA g4 (.ci(co0), .b(i21), .a(i11), .co(co), .o(o1));   //: @(561, 168) /sz:(130, 97) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Ro0<1 Ro1<1 ]
  //: input g3 (i22) @(164,296) /sn:0 /w:[ 1 ]
  //: input g2 (i21) @(163,264) /sn:0 /w:[ 0 ]
  //: input g1 (i12) @(163,184) /sn:0 /w:[ 0 ]
  //: output g6 (o1) @(853,214) /sn:0 /w:[ 0 ]
  //: output g7 (o2) @(855,259) /sn:0 /w:[ 1 ]
  HA g5 (.b(i22), .a(i12), .co(co0), .o(o2));   //: @(301, 299) /sz:(103, 90) /sn:0 /p:[ Li0>0 Li1>1 Ro0<0 Ro1<0 ]
  //: input g0 (i11) @(163,159) /sn:0 /w:[ 0 ]

endmodule
